.PARAM
+ LM1 = 4.653729365957649e-07
+ LM2 = 3.7079488855986813e-07
+ LM3 = 4.528365221742959e-07
+ LM4 = 4.6864854524782106e-07
+ LM5 = 2.3393927431056977e-07
+ LM6 = 4.762225257419609e-07
+ LM7 = 4.0727906188057457e-07
+ LM8 = 4.928810334270438e-07
+ WM1 = 5.402987794906587e-05
+ WM2 = 9.656709800221703e-06
+ WM3 = 3.0453596060637217e-05
+ WM4 = 2.5042732398990944e-05
+ WM5 = 4.2707455860015564e-05
+ WM6 = 3.6349845994253235e-05
+ WM7 = 4.46615864690664e-05
+ WM8 = 5.720284417026765e-05
