.PARAM
+ LM1 = 3.7355555317798267e-07
+ LM2 = 4.761214632100197e-07
+ LM3 = 4.984596182134089e-07
+ LM4 = 5.882044260865487e-07
+ LM5 = 3.094789855221767e-07
+ LM6 = 5.318561924269972e-07
+ LM7 = 5.38074396207641e-07
+ LM8 = 4.0504997339937196e-07
+ WM1 = 3.926766991025271e-05
+ WM2 = 4.057074273078096e-05
+ WM3 = 3.0054679847147e-05
+ WM4 = 5.282120337238513e-05
+ WM5 = 5.643256570540092e-05
+ WM6 = 4.554074354670248e-05
+ WM7 = 3.709223011379021e-05
+ WM8 = 4.9083236122342386e-05
