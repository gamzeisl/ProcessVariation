.PARAM
+ LM1 = 6.847709898678259e-07
+ LM2 = 8.5028125e-07
+ LM3 = 4.3346875e-07
+ WM1 = 5.179890625e-05
+ WM2 = 5.422015625e-05
+ WM3 = 9.42703125e-06
+ Ib = 0.00081746875
