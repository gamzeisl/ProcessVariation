.PARAM
+ LM1 = 2.558655060419944e-07
+ LM2 = 5.029810733360565e-07
+ LM3 = 2.0251211175225214e-07
+ LM4 = 6.337334789398807e-07
+ LM5 = 6.049902925327241e-07
+ LM6 = 4.142098986572279e-07
+ LM7 = 5.517775228590433e-07
+ LM8 = 3.3967994309319336e-07
+ WM1 = 4.977394444387989e-05
+ WM2 = 2.9327378940643162e-05
+ WM3 = 5.0067728421384144e-05
+ WM4 = 3.21823309625861e-05
+ WM5 = 1.880077856781465e-05
+ WM6 = 2.4861622090955936e-05
+ WM7 = 2.54901982494701e-05
+ WM8 = 2.201983147576424e-05
