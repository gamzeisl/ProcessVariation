.PARAM
+ LM1 = 5.82338108499601e-07
+ LM2 = 5.016636951665558e-07
+ LM3 = 4.045783268206528e-07
+ LM4 = 4.303007534684458e-07
+ LM5 = 2.7297700972736774e-07
+ LM6 = 4.499364704024497e-07
+ LM7 = 4.433467873640914e-07
+ LM8 = 2.014076204344522e-07
+ WM1 = 2.6871037102800586e-05
+ WM2 = 1.4107066930912307e-05
+ WM3 = 3.913995742187947e-05
+ WM4 = 2.205312616793194e-05
+ WM5 = 4.85398202602225e-05
+ WM6 = 3.2655644529840244e-05
+ WM7 = 6.234031102000232e-05
+ WM8 = 3.813303580838556e-05
