.PARAM
+ LM1 = 4.186568195518446e-07
+ LM2 = 4.844696109981899e-07
+ LM3 = 4.839230909408945e-07
+ LM4 = 5.804620199480064e-07
+ LM5 = 2.7897756814425854e-07
+ LM6 = 4.928132793380346e-07
+ LM7 = 5.626486540914132e-07
+ LM8 = 4.4063969975593876e-07
+ WM1 = 3.8422688051471476e-05
+ WM2 = 4.432321836779827e-05
+ WM3 = 3.305869179039813e-05
+ WM4 = 4.6420408116829366e-05
+ WM5 = 5.2040350663113445e-05
+ WM6 = 4.368046871624076e-05
+ WM7 = 2.609167780721404e-05
+ WM8 = 5.029650946541227e-05
