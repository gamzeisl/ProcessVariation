.PARAM
+ LM1 = 4.0881632197238813e-07
+ LM2 = 5.085711889740477e-07
+ LM3 = 3.854794762957038e-07
+ LM4 = 3.762606209568103e-07
+ LM5 = 5.811070162523021e-07
+ LM6 = 3.2997640092654346e-07
+ LM7 = 5.124995394970909e-07
+ LM8 = 3.8412552328267115e-07
+ WM1 = 5.128077999507378e-05
+ WM2 = 2.503262078622836e-05
+ WM3 = 5.149365677826501e-05
+ WM4 = 3.245844282667752e-05
+ WM5 = 2.5729284177540194e-05
+ WM6 = 4.442999738050951e-05
+ WM7 = 5.238462289950745e-05
+ WM8 = 9.471963042460188e-06
