.PARAM
+ LM1 = 4.873020672066172e-07
+ LM2 = 5.183661434562994e-07
+ LM3 = 5.735368233005245e-07
+ LM4 = 2.2720119618438363e-07
+ LM5 = 3.20596362351305e-07
+ LM6 = 4.760908489671529e-07
+ LM7 = 4.0555575031282544e-07
+ LM8 = 3.001141067798317e-07
+ WM1 = 3.334163200627185e-05
+ WM2 = 1.3864347973495079e-05
+ WM3 = 1.8959596037720023e-05
+ WM4 = 4.7648548434540635e-05
+ WM5 = 4.092636040253527e-05
+ WM6 = 2.7083387809792388e-05
+ WM7 = 6.014141237533121e-05
+ WM8 = 2.8845883569568533e-05
