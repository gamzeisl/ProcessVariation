.PARAM
+ LM1 = 1
+ LM2 = 2
+ LM3 = 3
+ LM4 = 4
+ LM5 = 5
+ LM6 = 6
