.PARAM
+ LM1 = 3.8359e-07
+ LM2 = 3.8379e-07
+ LM3 = 3.1352e-07
+ LM4 = 3.1353e-07
+ LM5 = 8.3656e-07
+ LM6 = 8.3594e-07
+ WM1 = 5.371e-05
+ WM2 = 5.3687e-05
+ WM3 = 7.4543e-05
+ WM4 = 7.455e-05
+ WM5 = 4.8142e-06
+ WM6 = 4.8145e-06
+ Rb = 2456.0316
+ Vb = 0.62019
