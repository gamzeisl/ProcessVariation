.PARAM
+ LM1 = 3.9426813777805473e-07
+ LM2 = 2.3232778663982204e-07
+ LM3 = 4.666652143503225e-07
+ LM4 = 4.5537556810045393e-07
+ LM5 = 2.3847225768356647e-07
+ LM6 = 6.087596044927942e-07
+ LM7 = 5.733862424835566e-07
+ LM8 = 4.2793282020234813e-07
+ WM1 = 3.305116397844902e-05
+ WM2 = 3.931665280914317e-05
+ WM3 = 4.538168205682013e-05
+ WM4 = 4.006357534321005e-05
+ WM5 = 5.759336957699168e-05
+ WM6 = 4.404642488127065e-05
+ WM7 = 4.9577851509003624e-05
+ WM8 = 9.900151279520014e-06
