.PARAM
+ LM1 = 5.141704856451022e-07
+ LM2 = 3.6376396124527395e-07
+ LM3 = 3.8408938089642277e-07
+ LM4 = 3.4931054854413685e-07
+ LM5 = 1.888133707443157e-07
+ LM6 = 5.121863372294543e-07
+ LM7 = 3.1723942030532215e-07
+ LM8 = 5.108013962376528e-07
+ WM1 = 5.561113270810613e-05
+ WM2 = 5.594766931420932e-05
+ WM3 = 1.592952099408997e-05
+ WM4 = 3.3697384519410046e-05
+ WM5 = 4.0317136246544016e-05
+ WM6 = 1.3349275857181318e-05
+ WM7 = 2.926966516484731e-05
+ WM8 = 6.024756407565162e-05
