.PARAM
+ LM1 = 1.0435187746357494e-06
+ LM2 = 7.749317737316132e-07
+ LM3 = 1.153167731256083e-06
+ WM1 = 5.095496694604118e-05
+ WM2 = 6.442705135453461e-05
+ WM3 = 7.214397107732786e-05
+ Ib = 0.0008029560114085484
