.PARAM
+ LM1 = 4.636177014524662e-07
+ LM2 = 4.510321663246159e-07
+ LM3 = 5.890585451829418e-07
+ LM4 = 2.3346989984238564e-07
+ LM5 = 3.119701743403547e-07
+ LM6 = 1.375458549714467e-07
+ LM7 = 4.380656140926917e-07
+ LM8 = 3.5674540672180566e-07
+ WM1 = 3.4886663725183956e-05
+ WM2 = 2.0166744443052792e-05
+ WM3 = 2.052002719645519e-05
+ WM4 = 1.8160545378371372e-05
+ WM5 = 3.5949084160658434e-05
+ WM6 = 2.993108289764999e-05
+ WM7 = 5.695079749758153e-05
+ WM8 = 2.1787662437352148e-05
