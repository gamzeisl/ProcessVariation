.PARAM
+ LM1 = 4.314336767372553e-07
+ LM2 = 4.2436368896567363e-07
+ LM3 = 3.9194165197013935e-07
+ LM4 = 4.123137002298834e-07
+ LM5 = 3.496100998665468e-07
+ LM6 = 4.4384608362960814e-07
+ LM7 = 4.0531475106725134e-07
+ LM8 = 5.167896539876418e-07
+ WM1 = 4.82559625179219e-05
+ WM2 = 8.869705710583862e-06
+ WM3 = 3.516187080289655e-05
+ WM4 = 3.640368264676672e-05
+ WM5 = 5.174172440260911e-05
+ WM6 = 2.3531613862163747e-05
+ WM7 = 2.7782331177765617e-05
+ WM8 = 5.280433477812846e-05
