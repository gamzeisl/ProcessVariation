.PARAM
+ LM1 = 1.09890625e-06
+ LM2 = 6.967187500000001e-07
+ LM3 = 7.3328125e-07
+ WM1 = 7.177421875e-05
+ WM2 = 2.334921875e-05
+ WM3 = 7.177421875e-05
+ Ib = 5.640625e-05
