.PARAM
+ LM1 = 3.525500457731098e-07
+ LM2 = 4.468149521664657e-07
+ LM3 = 4.3380638031031056e-07
+ LM4 = 4.771004575365025e-07
+ LM5 = 2.8310560427762065e-07
+ LM6 = 4.183987637417324e-07
+ LM7 = 4.965574498050914e-07
+ LM8 = 5.781594478912399e-07
+ WM1 = 4.3948658235599734e-05
+ WM2 = 1.0050475727372758e-05
+ WM3 = 4.4975105702287244e-05
+ WM4 = 2.8540797849236715e-05
+ WM5 = 3.654753859571996e-05
+ WM6 = 2.9877010920687252e-05
+ WM7 = 2.919224937764635e-05
+ WM8 = 4.8560167560729895e-05
