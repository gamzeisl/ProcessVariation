.PARAM
+ LM1 = 3.3478322416619123e-07
+ LM2 = 4.6184143267459474e-07
+ LM3 = 4.5680174005299935e-07
+ LM4 = 5.191375374660332e-07
+ LM5 = 2.654474713470486e-07
+ LM6 = 3.783256276227919e-07
+ LM7 = 5.358909255611319e-07
+ LM8 = 5.591219593333141e-07
+ WM1 = 2.104031305129291e-05
+ WM2 = 1.8913853891676358e-05
+ WM3 = 4.444931094916264e-05
+ WM4 = 3.104497921675237e-05
+ WM5 = 3.6622195160846044e-05
+ WM6 = 3.4914224634206505e-05
+ WM7 = 2.8769586035008453e-05
+ WM8 = 4.793321123255085e-05
