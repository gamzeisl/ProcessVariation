.PARAM
+ LM1 = 3.8401889991422955e-07
+ LM2 = 4.534320270753842e-07
+ LM3 = 5.038340424023627e-07
+ LM4 = 5.829072578253374e-07
+ LM5 = 4.013507270159177e-07
+ LM6 = 5.219279000458203e-07
+ LM7 = 5.263772263083655e-07
+ LM8 = 4.2264618002244103e-07
+ WM1 = 4.2152658718677605e-05
+ WM2 = 4.1880422222505614e-05
+ WM3 = 6.490983384074827e-06
+ WM4 = 4.9756796986198584e-05
+ WM5 = 5.389572362955168e-05
+ WM6 = 4.1811792734980575e-05
+ WM7 = 2.4261724415631438e-05
+ WM8 = 5.026151502996605e-05
