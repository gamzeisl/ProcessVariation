.PARAM
+ LM1 = 5.682159704307101e-07
+ LM2 = 2.9775592618635443e-07
+ LM3 = 2.804810984021749e-07
+ LM4 = 2.5119501761883396e-07
+ LM5 = 3.0672794951357293e-07
+ LM6 = 4.121763469717974e-07
+ LM7 = 4.970361119248604e-07
+ LM8 = 3.592759841603965e-07
+ WM1 = 4.8380455242419785e-05
+ WM2 = 5.0450166732501916e-05
+ WM3 = 1.121548405842938e-05
+ WM4 = 3.306637378214686e-05
+ WM5 = 2.947339696151207e-05
+ WM6 = 3.989604041128153e-05
+ WM7 = 3.913352824911027e-05
+ WM8 = 3.409690275373981e-05
