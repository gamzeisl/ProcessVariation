.PARAM
+ LM1 = 4.863794758088194e-07
+ LM2 = 3.3837541371597194e-07
+ LM3 = 7.352656154346933e-07
+ WM1 = 3.390615875090446e-05
+ WM2 = 9.325679925522646e-05
+ WM3 = 7.085096500017633e-05
+ Ib = 1.2040935341344074e-05
