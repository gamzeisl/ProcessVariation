.PARAM
+ LM1 = 4.7405574150122694e-07
+ LM2 = 4.897546467605078e-07
+ LM3 = 1.226424779185421e-06
+ WM1 = 9.245300389906665e-05
+ WM2 = 5.673204653563639e-05
+ WM3 = 4.946542846915434e-05
+ Ib = 0.0004906565577148835
