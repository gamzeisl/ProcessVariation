.PARAM
+ LM1 = 4.3116620313396176e-07
+ LM2 = 3.656179499887015e-07
+ LM3 = 1.9885445257516514e-07
+ LM4 = 4.919279683421983e-07
+ LM5 = 3.30696968228955e-07
+ LM6 = 5.566810243093929e-07
+ LM7 = 5.166243950389786e-07
+ LM8 = 5.581048390850597e-07
+ WM1 = 2.6804182370273677e-05
+ WM2 = 3.031392962281184e-05
+ WM3 = 3.874471568719578e-05
+ WM4 = 2.0558145212151452e-05
+ WM5 = 2.9157162086349407e-05
+ WM6 = 1.623391115769446e-05
+ WM7 = 3.802252613311476e-05
+ WM8 = 5.0020331405157066e-05
