.PARAM
+ LM1 = 5.890170574317451e-07
+ LM2 = 2.346436443397297e-07
+ LM3 = 2.214076593036582e-07
+ LM4 = 2.460054772163302e-07
+ LM5 = 4.615934196693375e-07
+ LM6 = 4.623469851438912e-07
+ LM7 = 6.223366979379656e-07
+ LM8 = 3.8078219862364376e-07
+ WM1 = 1.894978956069014e-05
+ WM2 = 5.9059274282624125e-05
+ WM3 = 2.6121192358227348e-05
+ WM4 = 5.237018453325562e-05
+ WM5 = 1.800954843636547e-05
+ WM6 = 2.537729633126704e-05
+ WM7 = 2.330515775732171e-05
+ WM8 = 3.5643726965919385e-05
