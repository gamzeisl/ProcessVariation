.PARAM
+ LM1 = 5.021354271430792e-07
+ LM2 = 6.720181387661821e-07
+ LM3 = 1.1669317055612677e-06
+ WM1 = 8.846890817996268e-05
+ WM2 = 6.198558489267494e-05
+ WM3 = 7.979814450913926e-06
+ Ib = 0.00024060750456985437
