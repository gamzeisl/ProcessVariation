.PARAM
+ LM1 = 4.698591044441388e-07
+ LM2 = 5.507657617103151e-07
+ LM3 = 8.674122281845475e-07
+ WM1 = 8.718057480522925e-05
+ WM2 = 3.161506959979167e-05
+ WM3 = 2.2242555020290854e-05
+ Ib = 0.0004727061118232755
